/*
 * Asynchronous FIFO with Gray Code Pointer Synchronization
 *
 * Implements a dual-clock FIFO for safe clock domain crossing.
 * Uses Gray code encoding for write/read pointers to ensure only
 * one bit changes at a time during synchronization.
 *
 * Features:
 *   - Independent write and read clock domains
 *   - Gray code pointer synchronization
 *   - Proper full/empty flag generation
 *   - Parameterizable width and depth (depth must be power of 2)
 *
 * Parameters:
 *   DATA_WIDTH - Width of data bus (default: 8)
 *   DEPTH      - FIFO depth, must be power of 2 (default: 8)
 *
 * Theory of Operation:
 *   - Write pointer increments in wr_clk domain
 *   - Read pointer increments in rd_clk domain
 *   - Pointers are converted to Gray code before synchronization
 *   - Only one bit changes in Gray code, safe for multi-bit CDC
 *   - Full flag generated by comparing synchronized rd_ptr in wr domain
 *   - Empty flag generated by comparing synchronized wr_ptr in rd domain
 */

module async_fifo #(
    parameter int DATA_WIDTH = 8,
    parameter int DEPTH = 8
) (
    // Write clock domain
    input  logic                    wr_clk,
    input  logic                    wr_rst_n,
    input  logic                    wr_clear,    // Synchronous clear in wr_clk domain
    input  logic                    wr_en,
    input  logic [DATA_WIDTH-1:0]   wr_data,
    output logic                    wr_full,
    output logic                    wr_almost_full,

    // Read clock domain
    input  logic                    rd_clk,
    input  logic                    rd_rst_n,
    input  logic                    rd_clear,    // Synchronous clear in rd_clk domain
    input  logic                    rd_en,
    output logic [DATA_WIDTH-1:0]   rd_data,
    output logic                    rd_empty,
    output logic                    rd_almost_empty
);

    // Calculate address width from depth
    localparam int ADDR_WIDTH = $clog2(DEPTH);
    localparam int PTR_WIDTH = ADDR_WIDTH + 1;  // Extra bit for full/empty detection

    // FIFO memory
    logic [DATA_WIDTH-1:0] mem [DEPTH-1:0];

    // Write domain pointers
    logic [PTR_WIDTH-1:0] wr_ptr;
    logic [PTR_WIDTH-1:0] wr_ptr_gray;
    logic [PTR_WIDTH-1:0] wr_ptr_gray_sync1;
    logic [PTR_WIDTH-1:0] wr_ptr_gray_sync2;

    // Read domain pointers
    logic [PTR_WIDTH-1:0] rd_ptr;
    logic [PTR_WIDTH-1:0] rd_ptr_gray;
    logic [PTR_WIDTH-1:0] rd_ptr_gray_sync1;
    logic [PTR_WIDTH-1:0] rd_ptr_gray_sync2;

    // Synchronized pointers (converted back to binary)
    logic [PTR_WIDTH-1:0] rd_ptr_sync;  // In write domain
    logic [PTR_WIDTH-1:0] wr_ptr_sync;  // In read domain

    //--------------------------------------------------------------------------
    // Binary to Gray Code Conversion
    //--------------------------------------------------------------------------

    function automatic logic [PTR_WIDTH-1:0] bin_to_gray(logic [PTR_WIDTH-1:0] bin);
        return bin ^ (bin >> 1);
    endfunction

    //--------------------------------------------------------------------------
    // Gray to Binary Code Conversion
    //--------------------------------------------------------------------------

    function automatic logic [PTR_WIDTH-1:0] gray_to_bin(logic [PTR_WIDTH-1:0] gray);
        logic [PTR_WIDTH-1:0] bin;
        bin[PTR_WIDTH-1] = gray[PTR_WIDTH-1];
        for (int i = PTR_WIDTH-2; i >= 0; i--) begin
            bin[i] = bin[i+1] ^ gray[i];
        end
        return bin;
    endfunction

    //--------------------------------------------------------------------------
    // Write Domain Logic
    //--------------------------------------------------------------------------

    // Write pointer and Gray code generation
    always_ff @(posedge wr_clk or negedge wr_rst_n) begin
        if (!wr_rst_n) begin
            wr_ptr <= '0;
            wr_ptr_gray <= '0;
        end else if (wr_clear) begin
            // Synchronous clear - reset pointers
            wr_ptr <= '0;
            wr_ptr_gray <= '0;
        end else if (wr_en && !wr_full) begin
            wr_ptr <= wr_ptr + 1'b1;
            wr_ptr_gray <= bin_to_gray(wr_ptr + 1'b1);
        end
    end

    // Synchronize read pointer to write domain (2-stage)
    always_ff @(posedge wr_clk or negedge wr_rst_n) begin
        if (!wr_rst_n) begin
            rd_ptr_gray_sync1 <= '0;
            rd_ptr_gray_sync2 <= '0;
        end else begin
            rd_ptr_gray_sync1 <= rd_ptr_gray;
            rd_ptr_gray_sync2 <= rd_ptr_gray_sync1;
        end
    end

    // Convert synchronized Gray read pointer back to binary
    assign rd_ptr_sync = gray_to_bin(rd_ptr_gray_sync2);

    // Full flag: write pointer has wrapped around and caught up to read pointer
    // Compare with extra MSB to distinguish full from empty
    assign wr_full = (wr_ptr[PTR_WIDTH-1] != rd_ptr_sync[PTR_WIDTH-1]) &&
                     (wr_ptr[PTR_WIDTH-2:0] == rd_ptr_sync[PTR_WIDTH-2:0]);

    // Almost full: one or two slots away from full
    logic [PTR_WIDTH-1:0] wr_ptr_next, wr_ptr_next2;
    assign wr_ptr_next = wr_ptr + {{(PTR_WIDTH-1){1'b0}}, 1'b1};
    assign wr_ptr_next2 = wr_ptr + {{(PTR_WIDTH-2){1'b0}}, 2'b10};

    assign wr_almost_full = ((wr_ptr_next[PTR_WIDTH-1] != rd_ptr_sync[PTR_WIDTH-1]) &&
                             (wr_ptr_next[PTR_WIDTH-2:0] == rd_ptr_sync[PTR_WIDTH-2:0])) ||
                            ((wr_ptr_next2[PTR_WIDTH-1] != rd_ptr_sync[PTR_WIDTH-1]) &&
                             (wr_ptr_next2[PTR_WIDTH-2:0] == rd_ptr_sync[PTR_WIDTH-2:0]));

    // Write to memory
    always_ff @(posedge wr_clk) begin
        if (wr_en && !wr_full) begin
            mem[wr_ptr[ADDR_WIDTH-1:0]] <= wr_data;
        end
    end

    //--------------------------------------------------------------------------
    // Read Domain Logic
    //--------------------------------------------------------------------------

    // Read pointer and Gray code generation
    always_ff @(posedge rd_clk or negedge rd_rst_n) begin
        if (!rd_rst_n) begin
            rd_ptr <= '0;
            rd_ptr_gray <= '0;
        end else if (rd_clear) begin
            // Synchronous clear - reset pointers
            rd_ptr <= '0;
            rd_ptr_gray <= '0;
        end else if (rd_en && !rd_empty) begin
            rd_ptr <= rd_ptr + 1'b1;
            rd_ptr_gray <= bin_to_gray(rd_ptr + 1'b1);
        end
    end

    // Synchronize write pointer to read domain (2-stage)
    always_ff @(posedge rd_clk or negedge rd_rst_n) begin
        if (!rd_rst_n) begin
            wr_ptr_gray_sync1 <= '0;
            wr_ptr_gray_sync2 <= '0;
        end else begin
            wr_ptr_gray_sync1 <= wr_ptr_gray;
            wr_ptr_gray_sync2 <= wr_ptr_gray_sync1;
        end
    end

    // Convert synchronized Gray write pointer back to binary
    assign wr_ptr_sync = gray_to_bin(wr_ptr_gray_sync2);

    // Empty flag: pointers are equal
    assign rd_empty = (rd_ptr == wr_ptr_sync);

    // Almost empty: one or two items left
    logic [PTR_WIDTH-1:0] rd_ptr_next, rd_ptr_next2;
    assign rd_ptr_next = rd_ptr + {{(PTR_WIDTH-1){1'b0}}, 1'b1};
    assign rd_ptr_next2 = rd_ptr + {{(PTR_WIDTH-2){1'b0}}, 2'b10};

    assign rd_almost_empty = (rd_ptr_next == wr_ptr_sync) ||
                             (rd_ptr_next2 == wr_ptr_sync);

    // Registered read output (standard FIFO behavior)
    // rd_data is valid one cycle after rd_en is asserted
    always_ff @(posedge rd_clk or negedge rd_rst_n) begin
        if (!rd_rst_n) begin
            rd_data <= '0;
        end else if (rd_en && !rd_empty) begin
            rd_data <= mem[rd_ptr[ADDR_WIDTH-1:0]];
        end
    end

    //--------------------------------------------------------------------------
    // Assertions
    //--------------------------------------------------------------------------

    // synthesis translate_off
    initial begin
        // Check that DEPTH is a power of 2
        assert ((DEPTH & (DEPTH - 1)) == 0) else
            $error("async_fifo: DEPTH must be a power of 2");

        assert (DEPTH >= 4) else
            $error("async_fifo: DEPTH must be at least 4");
    end

    // Check for overflow
    always @(posedge wr_clk) begin
        if (wr_rst_n && wr_en && wr_full) begin
            $error("async_fifo: Write to full FIFO!");
            $stop;
        end
    end

    // Check for underflow
    always @(posedge rd_clk) begin
        if (rd_rst_n && rd_en && rd_empty) begin
            $error("async_fifo: Read from empty FIFO!");
            $stop;
        end
    end
    // synthesis translate_on

endmodule
